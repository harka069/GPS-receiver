// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     Dec 15 2023 15:09:55

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    LED,
    clk,
    BUTTON3,
    BUTTON2,
    BUTTON1,
    BNC);

    output [9:0] LED;
    input clk;
    input BUTTON3;
    input BUTTON2;
    input BUTTON1;
    output BNC;

    wire N__1163;
    wire N__1162;
    wire N__1161;
    wire N__1152;
    wire N__1151;
    wire N__1150;
    wire N__1143;
    wire N__1142;
    wire N__1141;
    wire N__1134;
    wire N__1133;
    wire N__1132;
    wire N__1125;
    wire N__1124;
    wire N__1123;
    wire N__1116;
    wire N__1115;
    wire N__1114;
    wire N__1107;
    wire N__1106;
    wire N__1105;
    wire N__1098;
    wire N__1097;
    wire N__1096;
    wire N__1089;
    wire N__1088;
    wire N__1087;
    wire N__1080;
    wire N__1079;
    wire N__1078;
    wire N__1071;
    wire N__1070;
    wire N__1069;
    wire N__1062;
    wire N__1061;
    wire N__1060;
    wire N__1053;
    wire N__1052;
    wire N__1051;
    wire N__1044;
    wire N__1043;
    wire N__1042;
    wire N__1025;
    wire N__1024;
    wire N__1021;
    wire N__1018;
    wire N__1013;
    wire N__1010;
    wire N__1009;
    wire N__1006;
    wire N__1003;
    wire N__998;
    wire N__997;
    wire N__996;
    wire N__993;
    wire N__990;
    wire N__987;
    wire N__980;
    wire N__979;
    wire N__976;
    wire N__973;
    wire N__968;
    wire N__967;
    wire N__964;
    wire N__961;
    wire N__956;
    wire N__953;
    wire N__952;
    wire N__949;
    wire N__946;
    wire N__945;
    wire N__944;
    wire N__941;
    wire N__938;
    wire N__935;
    wire N__932;
    wire N__923;
    wire N__920;
    wire N__917;
    wire N__916;
    wire N__913;
    wire N__910;
    wire N__905;
    wire N__902;
    wire N__901;
    wire N__898;
    wire N__895;
    wire N__890;
    wire N__889;
    wire N__886;
    wire N__883;
    wire N__878;
    wire N__877;
    wire N__876;
    wire N__875;
    wire N__874;
    wire N__873;
    wire N__872;
    wire N__871;
    wire N__870;
    wire N__869;
    wire N__868;
    wire N__845;
    wire N__842;
    wire N__839;
    wire N__838;
    wire N__837;
    wire N__836;
    wire N__835;
    wire N__834;
    wire N__833;
    wire N__832;
    wire N__831;
    wire N__812;
    wire N__809;
    wire N__806;
    wire N__805;
    wire N__804;
    wire N__803;
    wire N__802;
    wire N__801;
    wire N__800;
    wire N__799;
    wire N__798;
    wire N__779;
    wire N__776;
    wire N__773;
    wire N__770;
    wire N__767;
    wire N__766;
    wire N__761;
    wire N__758;
    wire N__755;
    wire N__752;
    wire N__749;
    wire N__748;
    wire N__743;
    wire N__740;
    wire N__739;
    wire N__736;
    wire N__733;
    wire N__728;
    wire N__727;
    wire N__724;
    wire N__721;
    wire N__716;
    wire N__713;
    wire N__710;
    wire N__709;
    wire N__706;
    wire N__703;
    wire N__698;
    wire N__697;
    wire N__694;
    wire N__691;
    wire N__686;
    wire N__683;
    wire N__680;
    wire N__677;
    wire N__674;
    wire N__671;
    wire N__668;
    wire N__665;
    wire N__662;
    wire N__659;
    wire N__656;
    wire N__653;
    wire N__650;
    wire N__649;
    wire N__648;
    wire N__647;
    wire N__644;
    wire N__641;
    wire N__638;
    wire N__633;
    wire N__626;
    wire N__625;
    wire N__622;
    wire N__619;
    wire N__618;
    wire N__617;
    wire N__616;
    wire N__613;
    wire N__604;
    wire N__599;
    wire N__598;
    wire N__597;
    wire N__596;
    wire N__595;
    wire N__594;
    wire N__591;
    wire N__580;
    wire N__575;
    wire N__574;
    wire N__571;
    wire N__568;
    wire N__563;
    wire N__560;
    wire N__559;
    wire N__558;
    wire N__555;
    wire N__550;
    wire N__545;
    wire N__542;
    wire N__541;
    wire N__538;
    wire N__535;
    wire N__530;
    wire N__527;
    wire N__524;
    wire N__521;
    wire VCCG0;
    wire GNDG0;
    wire BUTTON1_c;
    wire BUTTON1_c_i;
    wire stevec_e_RNIL8L9Z0Z_4_cascade_;
    wire stevec_RNI8OFCZ0Z_1;
    wire LED_c_0;
    wire stevecZ0Z_2;
    wire stevecZ0Z_1;
    wire stevecZ0Z_0;
    wire stevec_i_4;
    wire stevecZ0Z_3;
    wire LED_c_1;
    wire \G2.qZ0Z_4 ;
    wire \G2.q_G2_2 ;
    wire \G2.q_G2_1 ;
    wire \G2.q_G2_5 ;
    wire \G2.q_G2_9 ;
    wire \G2.q_G2_8 ;
    wire \G2.data2_3 ;
    wire LED_c_3;
    wire q_G2_3;
    wire BUTTON3_c;
    wire BNC_c;
    wire \G2.q_G2_7 ;
    wire q_G2_6;
    wire LED_c_2;
    wire LED_c_5;
    wire LED_c_4;
    wire LED_c_9;
    wire LED_c_8;
    wire LED_c_7;
    wire LED_c_6;
    wire _gnd_net_;
    wire clk_0_c_g;
    wire N_31_g;
    wire BUTTON1_c_i_g;

    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__1161),
            .GLOBALBUFFEROUTPUT(clk_0_c_g));
    defparam clk_ibuf_gb_io_iopad.PULLUP=1'b0;
    defparam clk_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__1163),
            .DIN(N__1162),
            .DOUT(N__1161),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__1163),
            .PADOUT(N__1162),
            .PADIN(N__1161),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam BNC_obuf_iopad.PULLUP=1'b0;
    defparam BNC_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD BNC_obuf_iopad (
            .OE(N__1152),
            .DIN(N__1151),
            .DOUT(N__1150),
            .PACKAGEPIN(BNC));
    defparam BNC_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BNC_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BNC_obuf_preio (
            .PADOEN(N__1152),
            .PADOUT(N__1151),
            .PADIN(N__1150),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__677),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam BUTTON1_ibuf_iopad.PULLUP=1'b0;
    defparam BUTTON1_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD BUTTON1_ibuf_iopad (
            .OE(N__1143),
            .DIN(N__1142),
            .DOUT(N__1141),
            .PACKAGEPIN(BUTTON1));
    defparam BUTTON1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BUTTON1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BUTTON1_ibuf_preio (
            .PADOEN(N__1143),
            .PADOUT(N__1142),
            .PADIN(N__1141),
            .CLOCKENABLE(),
            .DIN0(BUTTON1_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam BUTTON3_ibuf_iopad.PULLUP=1'b0;
    defparam BUTTON3_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD BUTTON3_ibuf_iopad (
            .OE(N__1134),
            .DIN(N__1133),
            .DOUT(N__1132),
            .PACKAGEPIN(BUTTON3));
    defparam BUTTON3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BUTTON3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BUTTON3_ibuf_preio (
            .PADOEN(N__1134),
            .PADOUT(N__1133),
            .PADIN(N__1132),
            .CLOCKENABLE(),
            .DIN0(BUTTON3_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_obuf_0_iopad.PULLUP=1'b0;
    defparam LED_obuf_0_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED_obuf_0_iopad (
            .OE(N__1125),
            .DIN(N__1124),
            .DOUT(N__1123),
            .PACKAGEPIN(LED[0]));
    defparam LED_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam LED_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_obuf_0_preio (
            .PADOEN(N__1125),
            .PADOUT(N__1124),
            .PADIN(N__1123),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__656),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_obuf_1_iopad.PULLUP=1'b0;
    defparam LED_obuf_1_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED_obuf_1_iopad (
            .OE(N__1116),
            .DIN(N__1115),
            .DOUT(N__1114),
            .PACKAGEPIN(LED[1]));
    defparam LED_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam LED_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_obuf_1_preio (
            .PADOEN(N__1116),
            .PADOUT(N__1115),
            .PADIN(N__1114),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__545),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_obuf_2_iopad.PULLUP=1'b0;
    defparam LED_obuf_2_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED_obuf_2_iopad (
            .OE(N__1107),
            .DIN(N__1106),
            .DOUT(N__1105),
            .PACKAGEPIN(LED[2]));
    defparam LED_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam LED_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_obuf_2_preio (
            .PADOEN(N__1107),
            .PADOUT(N__1106),
            .PADIN(N__1105),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__998),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_obuf_3_iopad.PULLUP=1'b0;
    defparam LED_obuf_3_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED_obuf_3_iopad (
            .OE(N__1098),
            .DIN(N__1097),
            .DOUT(N__1096),
            .PACKAGEPIN(LED[3]));
    defparam LED_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam LED_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_obuf_3_preio (
            .PADOEN(N__1098),
            .PADOUT(N__1097),
            .PADIN(N__1096),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__710),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_obuf_4_iopad.PULLUP=1'b0;
    defparam LED_obuf_4_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED_obuf_4_iopad (
            .OE(N__1089),
            .DIN(N__1088),
            .DOUT(N__1087),
            .PACKAGEPIN(LED[4]));
    defparam LED_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam LED_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_obuf_4_preio (
            .PADOEN(N__1089),
            .PADOUT(N__1088),
            .PADIN(N__1087),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__968),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_obuf_5_iopad.PULLUP=1'b0;
    defparam LED_obuf_5_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED_obuf_5_iopad (
            .OE(N__1080),
            .DIN(N__1079),
            .DOUT(N__1078),
            .PACKAGEPIN(LED[5]));
    defparam LED_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam LED_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_obuf_5_preio (
            .PADOEN(N__1080),
            .PADOUT(N__1079),
            .PADIN(N__1078),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__980),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_obuf_6_iopad.PULLUP=1'b0;
    defparam LED_obuf_6_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED_obuf_6_iopad (
            .OE(N__1071),
            .DIN(N__1070),
            .DOUT(N__1069),
            .PACKAGEPIN(LED[6]));
    defparam LED_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam LED_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_obuf_6_preio (
            .PADOEN(N__1071),
            .PADOUT(N__1070),
            .PADIN(N__1069),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__890),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_obuf_7_iopad.PULLUP=1'b0;
    defparam LED_obuf_7_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED_obuf_7_iopad (
            .OE(N__1062),
            .DIN(N__1061),
            .DOUT(N__1060),
            .PACKAGEPIN(LED[7]));
    defparam LED_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam LED_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_obuf_7_preio (
            .PADOEN(N__1062),
            .PADOUT(N__1061),
            .PADIN(N__1060),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__905),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_obuf_8_iopad.PULLUP=1'b0;
    defparam LED_obuf_8_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED_obuf_8_iopad (
            .OE(N__1053),
            .DIN(N__1052),
            .DOUT(N__1051),
            .PACKAGEPIN(LED[8]));
    defparam LED_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam LED_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_obuf_8_preio (
            .PADOEN(N__1053),
            .PADOUT(N__1052),
            .PADIN(N__1051),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__923),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_obuf_9_iopad.PULLUP=1'b0;
    defparam LED_obuf_9_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED_obuf_9_iopad (
            .OE(N__1044),
            .DIN(N__1043),
            .DOUT(N__1042),
            .PACKAGEPIN(LED[9]));
    defparam LED_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam LED_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO LED_obuf_9_preio (
            .PADOEN(N__1044),
            .PADOUT(N__1043),
            .PADIN(N__1042),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__956),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__216 (
            .O(N__1025),
            .I(N__1021));
    InMux I__215 (
            .O(N__1024),
            .I(N__1018));
    LocalMux I__214 (
            .O(N__1021),
            .I(\G2.q_G2_7 ));
    LocalMux I__213 (
            .O(N__1018),
            .I(\G2.q_G2_7 ));
    CascadeMux I__212 (
            .O(N__1013),
            .I(N__1010));
    InMux I__211 (
            .O(N__1010),
            .I(N__1006));
    InMux I__210 (
            .O(N__1009),
            .I(N__1003));
    LocalMux I__209 (
            .O(N__1006),
            .I(q_G2_6));
    LocalMux I__208 (
            .O(N__1003),
            .I(q_G2_6));
    IoInMux I__207 (
            .O(N__998),
            .I(N__993));
    InMux I__206 (
            .O(N__997),
            .I(N__990));
    InMux I__205 (
            .O(N__996),
            .I(N__987));
    LocalMux I__204 (
            .O(N__993),
            .I(LED_c_2));
    LocalMux I__203 (
            .O(N__990),
            .I(LED_c_2));
    LocalMux I__202 (
            .O(N__987),
            .I(LED_c_2));
    IoInMux I__201 (
            .O(N__980),
            .I(N__976));
    InMux I__200 (
            .O(N__979),
            .I(N__973));
    LocalMux I__199 (
            .O(N__976),
            .I(LED_c_5));
    LocalMux I__198 (
            .O(N__973),
            .I(LED_c_5));
    IoInMux I__197 (
            .O(N__968),
            .I(N__964));
    InMux I__196 (
            .O(N__967),
            .I(N__961));
    LocalMux I__195 (
            .O(N__964),
            .I(LED_c_4));
    LocalMux I__194 (
            .O(N__961),
            .I(LED_c_4));
    IoInMux I__193 (
            .O(N__956),
            .I(N__953));
    LocalMux I__192 (
            .O(N__953),
            .I(N__949));
    InMux I__191 (
            .O(N__952),
            .I(N__946));
    Span4Mux_s2_h I__190 (
            .O(N__949),
            .I(N__941));
    LocalMux I__189 (
            .O(N__946),
            .I(N__938));
    InMux I__188 (
            .O(N__945),
            .I(N__935));
    InMux I__187 (
            .O(N__944),
            .I(N__932));
    Odrv4 I__186 (
            .O(N__941),
            .I(LED_c_9));
    Odrv4 I__185 (
            .O(N__938),
            .I(LED_c_9));
    LocalMux I__184 (
            .O(N__935),
            .I(LED_c_9));
    LocalMux I__183 (
            .O(N__932),
            .I(LED_c_9));
    IoInMux I__182 (
            .O(N__923),
            .I(N__920));
    LocalMux I__181 (
            .O(N__920),
            .I(N__917));
    IoSpan4Mux I__180 (
            .O(N__917),
            .I(N__913));
    InMux I__179 (
            .O(N__916),
            .I(N__910));
    Odrv4 I__178 (
            .O(N__913),
            .I(LED_c_8));
    LocalMux I__177 (
            .O(N__910),
            .I(LED_c_8));
    IoInMux I__176 (
            .O(N__905),
            .I(N__902));
    LocalMux I__175 (
            .O(N__902),
            .I(N__898));
    InMux I__174 (
            .O(N__901),
            .I(N__895));
    Odrv4 I__173 (
            .O(N__898),
            .I(LED_c_7));
    LocalMux I__172 (
            .O(N__895),
            .I(LED_c_7));
    IoInMux I__171 (
            .O(N__890),
            .I(N__886));
    InMux I__170 (
            .O(N__889),
            .I(N__883));
    LocalMux I__169 (
            .O(N__886),
            .I(LED_c_6));
    LocalMux I__168 (
            .O(N__883),
            .I(LED_c_6));
    ClkMux I__167 (
            .O(N__878),
            .I(N__845));
    ClkMux I__166 (
            .O(N__877),
            .I(N__845));
    ClkMux I__165 (
            .O(N__876),
            .I(N__845));
    ClkMux I__164 (
            .O(N__875),
            .I(N__845));
    ClkMux I__163 (
            .O(N__874),
            .I(N__845));
    ClkMux I__162 (
            .O(N__873),
            .I(N__845));
    ClkMux I__161 (
            .O(N__872),
            .I(N__845));
    ClkMux I__160 (
            .O(N__871),
            .I(N__845));
    ClkMux I__159 (
            .O(N__870),
            .I(N__845));
    ClkMux I__158 (
            .O(N__869),
            .I(N__845));
    ClkMux I__157 (
            .O(N__868),
            .I(N__845));
    GlobalMux I__156 (
            .O(N__845),
            .I(N__842));
    gio2CtrlBuf I__155 (
            .O(N__842),
            .I(clk_0_c_g));
    CEMux I__154 (
            .O(N__839),
            .I(N__812));
    CEMux I__153 (
            .O(N__838),
            .I(N__812));
    CEMux I__152 (
            .O(N__837),
            .I(N__812));
    CEMux I__151 (
            .O(N__836),
            .I(N__812));
    CEMux I__150 (
            .O(N__835),
            .I(N__812));
    CEMux I__149 (
            .O(N__834),
            .I(N__812));
    CEMux I__148 (
            .O(N__833),
            .I(N__812));
    CEMux I__147 (
            .O(N__832),
            .I(N__812));
    CEMux I__146 (
            .O(N__831),
            .I(N__812));
    GlobalMux I__145 (
            .O(N__812),
            .I(N__809));
    gio2CtrlBuf I__144 (
            .O(N__809),
            .I(N_31_g));
    SRMux I__143 (
            .O(N__806),
            .I(N__779));
    SRMux I__142 (
            .O(N__805),
            .I(N__779));
    SRMux I__141 (
            .O(N__804),
            .I(N__779));
    SRMux I__140 (
            .O(N__803),
            .I(N__779));
    SRMux I__139 (
            .O(N__802),
            .I(N__779));
    SRMux I__138 (
            .O(N__801),
            .I(N__779));
    SRMux I__137 (
            .O(N__800),
            .I(N__779));
    SRMux I__136 (
            .O(N__799),
            .I(N__779));
    SRMux I__135 (
            .O(N__798),
            .I(N__779));
    GlobalMux I__134 (
            .O(N__779),
            .I(N__776));
    gio2CtrlBuf I__133 (
            .O(N__776),
            .I(BUTTON1_c_i_g));
    InMux I__132 (
            .O(N__773),
            .I(N__770));
    LocalMux I__131 (
            .O(N__770),
            .I(\G2.qZ0Z_4 ));
    InMux I__130 (
            .O(N__767),
            .I(N__761));
    InMux I__129 (
            .O(N__766),
            .I(N__761));
    LocalMux I__128 (
            .O(N__761),
            .I(\G2.q_G2_2 ));
    InMux I__127 (
            .O(N__758),
            .I(N__755));
    LocalMux I__126 (
            .O(N__755),
            .I(\G2.q_G2_1 ));
    CascadeMux I__125 (
            .O(N__752),
            .I(N__749));
    InMux I__124 (
            .O(N__749),
            .I(N__743));
    InMux I__123 (
            .O(N__748),
            .I(N__743));
    LocalMux I__122 (
            .O(N__743),
            .I(\G2.q_G2_5 ));
    InMux I__121 (
            .O(N__740),
            .I(N__736));
    InMux I__120 (
            .O(N__739),
            .I(N__733));
    LocalMux I__119 (
            .O(N__736),
            .I(\G2.q_G2_9 ));
    LocalMux I__118 (
            .O(N__733),
            .I(\G2.q_G2_9 ));
    InMux I__117 (
            .O(N__728),
            .I(N__724));
    InMux I__116 (
            .O(N__727),
            .I(N__721));
    LocalMux I__115 (
            .O(N__724),
            .I(\G2.q_G2_8 ));
    LocalMux I__114 (
            .O(N__721),
            .I(\G2.q_G2_8 ));
    InMux I__113 (
            .O(N__716),
            .I(N__713));
    LocalMux I__112 (
            .O(N__713),
            .I(\G2.data2_3 ));
    IoInMux I__111 (
            .O(N__710),
            .I(N__706));
    InMux I__110 (
            .O(N__709),
            .I(N__703));
    LocalMux I__109 (
            .O(N__706),
            .I(LED_c_3));
    LocalMux I__108 (
            .O(N__703),
            .I(LED_c_3));
    InMux I__107 (
            .O(N__698),
            .I(N__694));
    InMux I__106 (
            .O(N__697),
            .I(N__691));
    LocalMux I__105 (
            .O(N__694),
            .I(q_G2_3));
    LocalMux I__104 (
            .O(N__691),
            .I(q_G2_3));
    InMux I__103 (
            .O(N__686),
            .I(N__683));
    LocalMux I__102 (
            .O(N__683),
            .I(N__680));
    Odrv12 I__101 (
            .O(N__680),
            .I(BUTTON3_c));
    IoInMux I__100 (
            .O(N__677),
            .I(N__674));
    LocalMux I__99 (
            .O(N__674),
            .I(N__671));
    Span4Mux_s2_h I__98 (
            .O(N__671),
            .I(N__668));
    Odrv4 I__97 (
            .O(N__668),
            .I(BNC_c));
    CascadeMux I__96 (
            .O(N__665),
            .I(stevec_e_RNIL8L9Z0Z_4_cascade_));
    IoInMux I__95 (
            .O(N__662),
            .I(N__659));
    LocalMux I__94 (
            .O(N__659),
            .I(stevec_RNI8OFCZ0Z_1));
    IoInMux I__93 (
            .O(N__656),
            .I(N__653));
    LocalMux I__92 (
            .O(N__653),
            .I(LED_c_0));
    CascadeMux I__91 (
            .O(N__650),
            .I(N__644));
    InMux I__90 (
            .O(N__649),
            .I(N__641));
    InMux I__89 (
            .O(N__648),
            .I(N__638));
    InMux I__88 (
            .O(N__647),
            .I(N__633));
    InMux I__87 (
            .O(N__644),
            .I(N__633));
    LocalMux I__86 (
            .O(N__641),
            .I(stevecZ0Z_2));
    LocalMux I__85 (
            .O(N__638),
            .I(stevecZ0Z_2));
    LocalMux I__84 (
            .O(N__633),
            .I(stevecZ0Z_2));
    CascadeMux I__83 (
            .O(N__626),
            .I(N__622));
    CascadeMux I__82 (
            .O(N__625),
            .I(N__619));
    InMux I__81 (
            .O(N__622),
            .I(N__613));
    InMux I__80 (
            .O(N__619),
            .I(N__604));
    InMux I__79 (
            .O(N__618),
            .I(N__604));
    InMux I__78 (
            .O(N__617),
            .I(N__604));
    InMux I__77 (
            .O(N__616),
            .I(N__604));
    LocalMux I__76 (
            .O(N__613),
            .I(stevecZ0Z_1));
    LocalMux I__75 (
            .O(N__604),
            .I(stevecZ0Z_1));
    InMux I__74 (
            .O(N__599),
            .I(N__591));
    InMux I__73 (
            .O(N__598),
            .I(N__580));
    InMux I__72 (
            .O(N__597),
            .I(N__580));
    InMux I__71 (
            .O(N__596),
            .I(N__580));
    InMux I__70 (
            .O(N__595),
            .I(N__580));
    InMux I__69 (
            .O(N__594),
            .I(N__580));
    LocalMux I__68 (
            .O(N__591),
            .I(stevecZ0Z_0));
    LocalMux I__67 (
            .O(N__580),
            .I(stevecZ0Z_0));
    InMux I__66 (
            .O(N__575),
            .I(N__571));
    InMux I__65 (
            .O(N__574),
            .I(N__568));
    LocalMux I__64 (
            .O(N__571),
            .I(stevec_i_4));
    LocalMux I__63 (
            .O(N__568),
            .I(stevec_i_4));
    CEMux I__62 (
            .O(N__563),
            .I(N__560));
    LocalMux I__61 (
            .O(N__560),
            .I(N__555));
    InMux I__60 (
            .O(N__559),
            .I(N__550));
    InMux I__59 (
            .O(N__558),
            .I(N__550));
    Odrv12 I__58 (
            .O(N__555),
            .I(stevecZ0Z_3));
    LocalMux I__57 (
            .O(N__550),
            .I(stevecZ0Z_3));
    IoInMux I__56 (
            .O(N__545),
            .I(N__542));
    LocalMux I__55 (
            .O(N__542),
            .I(N__538));
    InMux I__54 (
            .O(N__541),
            .I(N__535));
    Odrv4 I__53 (
            .O(N__538),
            .I(LED_c_1));
    LocalMux I__52 (
            .O(N__535),
            .I(LED_c_1));
    InMux I__51 (
            .O(N__530),
            .I(N__527));
    LocalMux I__50 (
            .O(N__527),
            .I(BUTTON1_c));
    IoInMux I__49 (
            .O(N__524),
            .I(N__521));
    LocalMux I__48 (
            .O(N__521),
            .I(BUTTON1_c_i));
    ICE_GB stevec_RNI8OFC_0_1 (
            .USERSIGNALTOGLOBALBUFFER(N__662),
            .GLOBALBUFFEROUTPUT(N_31_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB BUTTON1_ibuf_RNIIUI2_0 (
            .USERSIGNALTOGLOBALBUFFER(N__524),
            .GLOBALBUFFEROUTPUT(BUTTON1_c_i_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam BUTTON1_ibuf_RNIIUI2_LC_1_4_5.C_ON=1'b0;
    defparam BUTTON1_ibuf_RNIIUI2_LC_1_4_5.SEQ_MODE=4'b0000;
    defparam BUTTON1_ibuf_RNIIUI2_LC_1_4_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 BUTTON1_ibuf_RNIIUI2_LC_1_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__530),
            .lcout(BUTTON1_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam stevec_3_LC_1_5_0.C_ON=1'b0;
    defparam stevec_3_LC_1_5_0.SEQ_MODE=4'b1000;
    defparam stevec_3_LC_1_5_0.LUT_INIT=16'b0110101010101010;
    LogicCell40 stevec_3_LC_1_5_0 (
            .in0(N__559),
            .in1(N__648),
            .in2(N__625),
            .in3(N__598),
            .lcout(stevecZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__868),
            .ce(),
            .sr(_gnd_net_));
    defparam stevec_0_LC_1_5_2.C_ON=1'b0;
    defparam stevec_0_LC_1_5_2.SEQ_MODE=4'b1000;
    defparam stevec_0_LC_1_5_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 stevec_0_LC_1_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__596),
            .lcout(stevecZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__868),
            .ce(),
            .sr(_gnd_net_));
    defparam stevec_2_LC_1_5_3.C_ON=1'b0;
    defparam stevec_2_LC_1_5_3.SEQ_MODE=4'b1000;
    defparam stevec_2_LC_1_5_3.LUT_INIT=16'b0110011011001100;
    LogicCell40 stevec_2_LC_1_5_3 (
            .in0(N__595),
            .in1(N__647),
            .in2(_gnd_net_),
            .in3(N__618),
            .lcout(stevecZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__868),
            .ce(),
            .sr(_gnd_net_));
    defparam stevec_e_RNIL8L9_4_LC_1_5_4.C_ON=1'b0;
    defparam stevec_e_RNIL8L9_4_LC_1_5_4.SEQ_MODE=4'b0000;
    defparam stevec_e_RNIL8L9_4_LC_1_5_4.LUT_INIT=16'b0000000010000000;
    LogicCell40 stevec_e_RNIL8L9_4_LC_1_5_4 (
            .in0(N__558),
            .in1(N__594),
            .in2(N__650),
            .in3(N__574),
            .lcout(),
            .ltout(stevec_e_RNIL8L9Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam stevec_RNI8OFC_1_LC_1_5_5.C_ON=1'b0;
    defparam stevec_RNI8OFC_1_LC_1_5_5.SEQ_MODE=4'b0000;
    defparam stevec_RNI8OFC_1_LC_1_5_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 stevec_RNI8OFC_1_LC_1_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__665),
            .in3(N__616),
            .lcout(stevec_RNI8OFCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam stevec_1_LC_1_5_6.C_ON=1'b0;
    defparam stevec_1_LC_1_5_6.SEQ_MODE=4'b1000;
    defparam stevec_1_LC_1_5_6.LUT_INIT=16'b0101010110101010;
    LogicCell40 stevec_1_LC_1_5_6 (
            .in0(N__617),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__597),
            .lcout(stevecZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__868),
            .ce(),
            .sr(_gnd_net_));
    defparam \G1.q_0_LC_1_7_5 .C_ON=1'b0;
    defparam \G1.q_0_LC_1_7_5 .SEQ_MODE=4'b1011;
    defparam \G1.q_0_LC_1_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G1.q_0_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__541),
            .lcout(LED_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__870),
            .ce(N__832),
            .sr(N__798));
    defparam stevec_e_4_LC_2_5_0.C_ON=1'b0;
    defparam stevec_e_4_LC_2_5_0.SEQ_MODE=4'b1000;
    defparam stevec_e_4_LC_2_5_0.LUT_INIT=16'b0110101010101010;
    LogicCell40 stevec_e_4_LC_2_5_0 (
            .in0(N__575),
            .in1(N__649),
            .in2(N__626),
            .in3(N__599),
            .lcout(stevec_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__869),
            .ce(N__563),
            .sr(_gnd_net_));
    defparam \G1.q_1_LC_2_7_5 .C_ON=1'b0;
    defparam \G1.q_1_LC_2_7_5 .SEQ_MODE=4'b1011;
    defparam \G1.q_1_LC_2_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G1.q_1_LC_2_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__997),
            .lcout(LED_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__872),
            .ce(N__833),
            .sr(N__800));
    defparam \G2.q_8_LC_3_5_0 .C_ON=1'b0;
    defparam \G2.q_8_LC_3_5_0 .SEQ_MODE=4'b1011;
    defparam \G2.q_8_LC_3_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G2.q_8_LC_3_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__740),
            .lcout(\G2.q_G2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__871),
            .ce(N__831),
            .sr(N__799));
    defparam \G2.q_2_LC_3_5_1 .C_ON=1'b0;
    defparam \G2.q_2_LC_3_5_1 .SEQ_MODE=4'b1011;
    defparam \G2.q_2_LC_3_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G2.q_2_LC_3_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__697),
            .lcout(\G2.q_G2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__871),
            .ce(N__831),
            .sr(N__799));
    defparam \G2.q_4_LC_3_5_2 .C_ON=1'b0;
    defparam \G2.q_4_LC_3_5_2 .SEQ_MODE=4'b1011;
    defparam \G2.q_4_LC_3_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G2.q_4_LC_3_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__748),
            .lcout(\G2.qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__871),
            .ce(N__831),
            .sr(N__799));
    defparam \G2.q_7_LC_3_5_3 .C_ON=1'b0;
    defparam \G2.q_7_LC_3_5_3 .SEQ_MODE=4'b1011;
    defparam \G2.q_7_LC_3_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G2.q_7_LC_3_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__728),
            .lcout(\G2.q_G2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__871),
            .ce(N__831),
            .sr(N__799));
    defparam \G2.q_5_LC_3_5_4 .C_ON=1'b0;
    defparam \G2.q_5_LC_3_5_4 .SEQ_MODE=4'b1011;
    defparam \G2.q_5_LC_3_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G2.q_5_LC_3_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1009),
            .lcout(\G2.q_G2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__871),
            .ce(N__831),
            .sr(N__799));
    defparam \G2.q_3_LC_3_5_5 .C_ON=1'b0;
    defparam \G2.q_3_LC_3_5_5 .SEQ_MODE=4'b1011;
    defparam \G2.q_3_LC_3_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G2.q_3_LC_3_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__773),
            .lcout(q_G2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__871),
            .ce(N__831),
            .sr(N__799));
    defparam \G2.q_1_LC_3_5_6 .C_ON=1'b0;
    defparam \G2.q_1_LC_3_5_6 .SEQ_MODE=4'b1011;
    defparam \G2.q_1_LC_3_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G2.q_1_LC_3_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__767),
            .lcout(\G2.q_G2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__871),
            .ce(N__831),
            .sr(N__799));
    defparam \G2.q_9_LC_3_5_7 .C_ON=1'b0;
    defparam \G2.q_9_LC_3_5_7 .SEQ_MODE=4'b1011;
    defparam \G2.q_9_LC_3_5_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \G2.q_9_LC_3_5_7  (
            .in0(N__766),
            .in1(N__758),
            .in2(N__752),
            .in3(N__716),
            .lcout(\G2.q_G2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__871),
            .ce(N__831),
            .sr(N__799));
    defparam \G2.q_RNO_0_9_LC_3_6_3 .C_ON=1'b0;
    defparam \G2.q_RNO_0_9_LC_3_6_3 .SEQ_MODE=4'b0000;
    defparam \G2.q_RNO_0_9_LC_3_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \G2.q_RNO_0_9_LC_3_6_3  (
            .in0(N__739),
            .in1(N__727),
            .in2(_gnd_net_),
            .in3(N__1024),
            .lcout(\G2.data2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \G1.q_2_LC_3_8_0 .C_ON=1'b0;
    defparam \G1.q_2_LC_3_8_0 .SEQ_MODE=4'b1011;
    defparam \G1.q_2_LC_3_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G1.q_2_LC_3_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__709),
            .lcout(LED_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__874),
            .ce(N__835),
            .sr(N__802));
    defparam \G1.q_3_LC_3_8_2 .C_ON=1'b0;
    defparam \G1.q_3_LC_3_8_2 .SEQ_MODE=4'b1011;
    defparam \G1.q_3_LC_3_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G1.q_3_LC_3_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__967),
            .lcout(LED_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__874),
            .ce(N__835),
            .sr(N__802));
    defparam BNC_obuf_RNO_LC_4_5_6.C_ON=1'b0;
    defparam BNC_obuf_RNO_LC_4_5_6.SEQ_MODE=4'b0000;
    defparam BNC_obuf_RNO_LC_4_5_6.LUT_INIT=16'b1110110100010010;
    LogicCell40 BNC_obuf_RNO_LC_4_5_6 (
            .in0(N__698),
            .in1(N__686),
            .in2(N__1013),
            .in3(N__952),
            .lcout(BNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \G2.q_6_LC_4_6_0 .C_ON=1'b0;
    defparam \G2.q_6_LC_4_6_0 .SEQ_MODE=4'b1011;
    defparam \G2.q_6_LC_4_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G2.q_6_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1025),
            .lcout(q_G2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__873),
            .ce(N__834),
            .sr(N__801));
    defparam \G1.q_9_LC_4_7_3 .C_ON=1'b0;
    defparam \G1.q_9_LC_4_7_3 .SEQ_MODE=4'b1011;
    defparam \G1.q_9_LC_4_7_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \G1.q_9_LC_4_7_3  (
            .in0(_gnd_net_),
            .in1(N__944),
            .in2(_gnd_net_),
            .in3(N__996),
            .lcout(LED_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__875),
            .ce(N__836),
            .sr(N__803));
    defparam \G1.q_5_LC_4_8_1 .C_ON=1'b0;
    defparam \G1.q_5_LC_4_8_1 .SEQ_MODE=4'b1011;
    defparam \G1.q_5_LC_4_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G1.q_5_LC_4_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__889),
            .lcout(LED_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__876),
            .ce(N__837),
            .sr(N__804));
    defparam \G1.q_4_LC_4_8_6 .C_ON=1'b0;
    defparam \G1.q_4_LC_4_8_6 .SEQ_MODE=4'b1011;
    defparam \G1.q_4_LC_4_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G1.q_4_LC_4_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__979),
            .lcout(LED_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__876),
            .ce(N__837),
            .sr(N__804));
    defparam \G1.q_7_LC_5_7_5 .C_ON=1'b0;
    defparam \G1.q_7_LC_5_7_5 .SEQ_MODE=4'b1011;
    defparam \G1.q_7_LC_5_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G1.q_7_LC_5_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__916),
            .lcout(LED_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__877),
            .ce(N__838),
            .sr(N__805));
    defparam \G1.q_8_LC_5_7_6 .C_ON=1'b0;
    defparam \G1.q_8_LC_5_7_6 .SEQ_MODE=4'b1011;
    defparam \G1.q_8_LC_5_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G1.q_8_LC_5_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__945),
            .lcout(LED_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__877),
            .ce(N__838),
            .sr(N__805));
    defparam \G1.q_6_LC_5_8_6 .C_ON=1'b0;
    defparam \G1.q_6_LC_5_8_6 .SEQ_MODE=4'b1011;
    defparam \G1.q_6_LC_5_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \G1.q_6_LC_5_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__901),
            .lcout(LED_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__878),
            .ce(N__839),
            .sr(N__806));
endmodule // TOP
